module Control_Unit(input [1:0] mode, input [3:0] OPCode, input S);

endmodule