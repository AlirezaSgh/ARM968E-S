module test(input PIN_N25, output PIN_AE23);
assign PIN_AE23 = PIN_N25;
endmodule
